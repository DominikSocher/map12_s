--------------------------------------------------
-- Inverter
-------------------------------------------------
library ieee;
use ieee.std_logic_1164.all; 

entity inv_a is
    port (
        i : in  std_logic;
        q : out std_logic     
    );
end entity inv_a;

architecture rtl of inv_a is
    
begin
    
    
    
end architecture rtl;