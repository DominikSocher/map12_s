--------------------------------------------------
-- or gate
-------------------------------------------------
library ieee;
use ieee.std_logic_1164.all; 

entity or_4 is
    port (
        i0 : in  std_logic;
        i1 : in  std_logic;
        i2 : in  std_logic;
        i3 : in  std_logic;
        q  : out std_logic         
    );
end entity or_4;

architecture rtl of or_4 is
    
begin
    
    
    
end architecture rtl;